`default_nettype none
module hart #(
    // After reset, the program counter (PC) should be initialized to this
    // address and start executing instructions from there.
    parameter RESET_ADDR = 32'h00000000
) (
    // Global clock.
    input  wire        i_clk,
    // Synchronous active-high reset.
    input  wire        i_rst,
    // Instruction fetch goes through a read only instruction memory (imem)
    // port. The port accepts a 32-bit address (e.g. from the program counter)
    // per cycle and combinationally returns a 32-bit instruction word. This
    // is not representative of a realistic memory interface; it has been
    // modeled as more similar to a DFF or SRAM to simplify phase 3. In
    // later phases, you will replace this with a more realistic memory.
    //
    // 32-bit read address for the instruction memory. This is expected to be
    // 4 byte aligned - that is, the two LSBs should be zero.
    output wire [31:0] o_imem_raddr,
    // Instruction word fetched from memory, available synchronously after
    // the next clock edge.
    // NOTE: This is different from the previous phase. To accomodate a
    // multi-cycle pipelined design, the instruction memory read is
    // now synchronous.
    input  wire [31:0] i_imem_rdata,
    // Data memory accesses go through a separate read/write data memory (dmem)
    // that is shared between read (load) and write (stored). The port accepts
    // a 32-bit address, read or write enable, and mask (explained below) each
    // cycle. Reads are combinational - values are available immediately after
    // updating the address and asserting read enable. Writes occur on (and
    // are visible at) the next clock edge.
    //
    // Read/write address for the data memory. This should be 32-bit aligned
    // (i.e. the two LSB should be zero). See `o_dmem_mask` for how to perform
    // half-word and byte accesses at unaligned addresses.
    output wire [31:0] o_dmem_addr,
    // When asserted, the memory will perform a read at the aligned address
    // specified by `i_addr` and return the 32-bit word at that address
    // immediately (i.e. combinationally). It is illegal to assert this and
    // `o_dmem_wen` on the same cycle.
    output wire        o_dmem_ren,
    // When asserted, the memory will perform a write to the aligned address
    // `o_dmem_addr`. When asserted, the memory will write the bytes in
    // `o_dmem_wdata` (specified by the mask) to memory at the specified
    // address on the next rising clock edge. It is illegal to assert this and
    // `o_dmem_ren` on the same cycle.
    output wire        o_dmem_wen,
    // The 32-bit word to write to memory when `o_dmem_wen` is asserted. When
    // write enable is asserted, the byte lanes specified by the mask will be
    // written to the memory word at the aligned address at the next rising
    // clock edge. The other byte lanes of the word will be unaffected.
    output wire [31:0] o_dmem_wdata,
    // The dmem interface expects word (32 bit) aligned addresses. However,
    // WISC-25 supports byte and half-word loads and stores at unaligned and
    // 16-bit aligned addresses, respectively. To support this, the access
    // mask specifies which bytes within the 32-bit word are actually read
    // from or written to memory.
    //
    // To perform a half-word read at address 0x00001002, align `o_dmem_addr`
    // to 0x00001000, assert `o_dmem_ren`, and set the mask to 0b1100 to
    // indicate that only the upper two bytes should be read. Only the upper
    // two bytes of `i_dmem_rdata` can be assumed to have valid data; to
    // calculate the final value of the `lh[u]` instruction, shift the rdata
    // word right by 16 bits and sign/zero extend as appropriate.
    //
    // To perform a byte write at address 0x00002003, align `o_dmem_addr` to
    // `0x00002000`, assert `o_dmem_wen`, and set the mask to 0b1000 to
    // indicate that only the upper byte should be written. On the next clock
    // cycle, the upper byte of `o_dmem_wdata` will be written to memory, with
    // the other three bytes of the aligned word unaffected. Remember to shift
    // the value of the `sb` instruction left by 24 bits to place it in the
    // appropriate byte lane.
    output wire [ 3:0] o_dmem_mask,
    // The 32-bit word read from data memory. When `o_dmem_ren` is asserted,
    // after the next clock edge, this will reflect the contents of memory
    // at the specified address, for the bytes enabled by the mask. When
    // read enable is not asserted, or for bytes not set in the mask, the
    // value is undefined.
    // NOTE: This is different from the previous phase. To accomodate a
    // multi-cycle pipelined design, the data memory read is
    // now synchronous.
    input  wire [31:0] i_dmem_rdata,
	// The output `retire` interface is used to signal to the testbench that
    // the CPU has completed and retired an instruction. A single cycle
    // implementation will assert this every cycle; however, a pipelined
    // implementation that needs to stall (due to internal hazards or waiting
    // on memory accesses) will not assert the signal on cycles where the
    // instruction in the writeback stage is not retiring.
    //
    // Asserted when an instruction is being retired this cycle. If this is
    // not asserted, the other retire signals are ignored and may be left invalid.
    output wire        o_retire_valid,
    // The 32 bit instruction word of the instrution being retired. This
    // should be the unmodified instruction word fetched from instruction
    // memory.
    output wire [31:0] o_retire_inst,
    // Asserted if the instruction produced a trap, due to an illegal
    // instruction, unaligned data memory access, or unaligned instruction
    // address on a taken branch or jump.
    output wire        o_retire_trap,
    // Asserted if the instruction is an `ebreak` instruction used to halt the
    // processor. This is used for debugging and testing purposes to end
    // a program.
    output wire        o_retire_halt,
    // The first register address read by the instruction being retired. If
    // the instruction does not read from a register (like `lui`), this
    // should be 5'd0.
    output wire [ 4:0] o_retire_rs1_raddr,
    // The second register address read by the instruction being retired. If
    // the instruction does not read from a second register (like `addi`), this
    // should be 5'd0.
    output wire [ 4:0] o_retire_rs2_raddr,
    // The first source register data read from the register file (in the
    // decode stage) for the instruction being retired. If rs1 is 5'd0, this
    // should also be 32'd0.
    output wire [31:0] o_retire_rs1_rdata,
    // The second source register data read from the register file (in the
    // decode stage) for the instruction being retired. If rs2 is 5'd0, this
    // should also be 32'd0.
    output wire [31:0] o_retire_rs2_rdata,
    // The destination register address written by the instruction being
    // retired. If the instruction does not write to a register (like `sw`),
    // this should be 5'd0.
    output wire [ 4:0] o_retire_rd_waddr,
    // The destination register data written to the register file in the
    // writeback stage by this instruction. If rd is 5'd0, this field is
    // ignored and can be treated as a don't care.
    output wire [31:0] o_retire_rd_wdata,
    // The following data memory retire interface is used to record the
    // memory transactions completed by the instruction being retired.
    // As such, it mirrors the transactions happening on the main data
    // memory interface (o_dmem_* and i_dmem_*) but is delayed to match
    // the retirement of the instruction. You can hook this up by just
    // registering the main dmem interface signals into the writeback
    // stage of your pipeline.
    //
    // All these fields are don't-care for instructions that do not
    // access data memory (o_retire_dmem_ren and o_retire_dmem_wen
    // not asserted).
    // NOTE: This interface is new for phase 5 in order to account for
    // the delay between data memory accesses and instruction retire.
    //
    // The 32-bit data memory address accessed by the instruction.
    output wire [31:0] o_retire_dmem_addr,
    // The byte masked used for the data memory access.
    output wire [ 3:0] o_retire_dmem_mask,
    // Asserted if the instruction performed a read (load) from data memory.
    output wire        o_retire_dmem_ren,
    // Asserted if the instruction performed a write (store) to data memory.
    output wire        o_retire_dmem_wen,
    // The 32-bit data read from memory by a load instruction.
    output wire [31:0] o_retire_dmem_rdata,
    // The 32-bit data written to memory by a store instruction.
    output wire [31:0] o_retire_dmem_wdata,
    // The current program counter of the instruction being retired - i.e.
    // the instruction memory address that the instruction was fetched from.
    output wire [31:0] o_retire_pc,
    // the next program counter after the instruction is retired. For most
    // instructions, this is `o_retire_pc + 4`, but must be the branch or jump
    // target for *taken* branches and jumps.
    output wire [31:0] o_retire_next_pc

`ifdef RISCV_FORMAL
    ,`RVFI_OUTPUTS,
`endif
);


  /*
Delcleration of any extra wires needed for connecting modules and for signals used across modules 
*/

  wire [31:0] JB_PC;
  wire [31:0] current_PC;  //will hold current PC value 
  wire [31:0] next_PC;  //holds the adress to be updated in PC next 
  wire [31:0] PC_plus4;  //will hold PC+4 value

  wire        jal_C;  //control signal 
  wire        jalr_C;  //control signal 
  wire        branch_C;  //control signal 
  wire        MemRead_C;  //control signal 
  wire        MemWrite_C;  //control signal 
  wire [ 1:0] Data_sel_C;  //control signal 
  wire [ 2:0] ALUop_C;  //control signal 
  wire [31:0] ALU_operand1;  //alu operand 1
  wire [31:0] ALU_operand2;  //alu operand 2
  wire [31:0] immediate_val;  //generated immeidate 
  wire [31:0] Mem_WD;  //feeds into memory write data port 
  wire [ 2:0] func3_val;  //feeds into branch logic block
  wire [ 3:0] func_val;  //feeds into ALU control block

  wire [31:0] ALU_result;  //ALU operation result
  wire [ 1:0] PC_MUX_SEL;  //MUX select signal for choosing next PC
  wire [31:0] PC_offset;  //PC + immediate offset value
  wire [31:0] MEM_DATA;  //Data returned from memory read  
  wire [31:0] WB_DATA;  //data to be input into register file 
  wire IF_ID_En;  

  reg reg2_regWrite;
  reg [31:0] reg3_curr_instruct;

  /* 
 Instantiate IF section of proccesor 
*/


  // choose between PC+4 or jump/Branch PC (By default should be PC+4)
  reg rst_reg;
  assign next_PC =(rst_reg)?(32'd0):((~IF_ID_En)?(PC_plus4-32'd4):((PC_MUX_SEL[0]) ? JB_PC : PC_plus4));


  wire[31:0] current_PC_w;
  IF fetch_inst (
      .IF_EN(IF_ID_En),
      .i_clk   (i_clk),   //input- clk to control PC update
      .i_rst   (i_rst),   //input- used to reset PC to starting value
      .i_NextPC(next_PC), //input- next PC value                           

      .o_PC(current_PC_w),            //output- current PC feed into instruction memory and other locations (schematic) 
      .o_inc_pc(PC_plus4)  //output- current PC + 4 
  );
  assign current_PC=(IF_ID_En)?(current_PC_w):(current_PC_w-32'd4);

  assign o_imem_raddr = next_PC;  //assign instruction memory read adress to current PC


  /* 
 IF/ID Piepline Register
 Include NOP control
 TODO: EXPECTS INPUT OF NOP
*/
  reg[31:0] PC_plus4_flop;
  always@(posedge i_clk)begin
    if(i_rst)
      rst_reg<=1'b1;
    else
      rst_reg<=1'b0;
  end

reg [31:0] flopped_current_PC;
  always @(posedge i_clk) begin
    if (i_rst || rst_reg)begin
      flopped_current_PC      <= 32'd0;
    PC_plus4_flop<=32'd0;
  end
  else if (IF_ID_En)begin
      flopped_current_PC      <= current_PC;
    PC_plus4_flop<=PC_plus4;
  end
  else begin
      flopped_current_PC      <= flopped_current_PC; 
      PC_plus4_flop<=PC_plus4_flop;
    end
  end

  wire flush;
  //TODO: 
  reg reg1_jal_C;
  reg reg0_jal_C;
  reg reg0_jalr_C;
  assign flush=(reg0_jal_C ||reg0_jalr_C);

  reg [31:0] reg0_PC_plus4;
  reg [31:0] reg0_current_PC;
  reg [31:0] reg0_curr_instruct;

  reg reg0_retire_valid; 
  always @(posedge i_clk) begin
    if (i_rst || rst_reg||flush) begin
      reg0_PC_plus4      <= 32'd0;
      reg0_current_PC    <= 32'd0;
      reg0_curr_instruct <= 32'd0;
      reg0_retire_valid  <= 1'd0; 
    end else if (IF_ID_En) begin
      reg0_PC_plus4      <= PC_plus4;
      reg0_current_PC    <= current_PC;
      reg0_curr_instruct <= i_imem_rdata;
      reg0_retire_valid  <= 1'd1;
    end else begin 
      reg0_PC_plus4      <= reg0_PC_plus4;
      reg0_current_PC    <= reg0_current_PC;
      reg0_curr_instruct <= reg0_curr_instruct;
      reg0_retire_valid  <= reg0_retire_valid; 
    end
  end
  wire [4:0] IF_ID_RS1;
  wire [4:0] IF_ID_RS2;

  //input
  wire [4:0] ID_EX_WriteReg;
  wire ID_EX_RegWrite;

  wire [4:0] EX_MEM_WriteReg;
  wire EX_MEM_RegWrite;
  reg reg0_regWrite;
  reg [31:0] reg1_curr_instruct;
  reg [31:0] reg2_curr_instruct;
  reg reg1_regWrite; 

  //output
  wire PC_En;
  wire Mux_sel;
  //NOTE: diagram does NOT show this?
  hazard haz (
  .op_code(reg0_curr_instruct[6:0]),
      .IF_ID_RS1(reg0_curr_instruct[19:15]),
      .IF_ID_RS2(reg0_curr_instruct[24:20]),
      .ID_EX_RegWrite(reg0_regWrite),
      .EX_MEM_RegWrite(reg1_regWrite), 
      .ID_EX_WriteReg(reg1_curr_instruct[11:7]),
      .EX_MEM_WriteReg(reg2_curr_instruct[11:7]),
      .valid_inst(reg0_retire_valid),

      .PC_En(PC_En),
      .IF_ID_En(IF_ID_En),
      .Mux_sel(Mux_sel)
  );

  /* 
 Instantiate ID section of proccesor 
*/

  //////////Internal Wires////////////
  //to connect top-level register file to decode block
  wire [31:0] regData1;
  wire [31:0] regData2;
  wire regWrite;

  ID decode_I (
      .rst        (i_rst),               //input- to RF
      .clk        (i_clk),               //input- to RF
      .i_instruct (reg0_curr_instruct),  //input- full instruction input
      .i_currentPC(reg0_current_PC),     //input- the current PC value (used for auipc instruction)
      .o_RegWrite (regWrite),
      .i_regData1 (regData1),
      .i_regData2 (regData2),
      .o_jal     (jal_C),          //output- from control unit
      .o_jalr    (jalr_C),         //output- from control unit
      .o_branch  (branch_C),       //output- from control unit
      .o_MemRead (MemRead_C),      //output- from control unit
      .o_Data_sel(Data_sel_C),     //output- from control unit used for WB module
      .o_MemWrite(MemWrite_C),     //output- from control unit
      .o_op1     (ALU_operand1),   //output- from control unit (select ALU operand)
      .o_op2     (ALU_operand2),   //output- from control unit (selects ALU operand)
      .o_ALUop   (ALUop_C),        //output- from control unit goes to ALU control
      .o_imm     (immediate_val),  //output- the generated immediate 
      .o_Rdata2  (Mem_WD),         //output- will feed into memory 'write data' port 
      .func      (func_val),       //output- combination of func7 and func3 for ALU control block
      .func3     (func3_val)       //output- func 3 for branch logic 
  );

  //write adress should be 0 when instruction does not write to register 
  wire [4:0] rf_writeAddress;
  assign rf_writeAddress = (reg2_regWrite) ? reg3_curr_instruct[11:7] : 5'b00000;

  wire [31:0] WriteDataReg;
  rf rf (
      .i_clk(i_clk),
      .i_rst(i_rst),

      .i_rs1_raddr(reg0_curr_instruct[19:15]),
      .i_rs2_raddr(reg0_curr_instruct[24:20]),

      .o_rs1_rdata(regData1),
      .o_rs2_rdata(regData2),

      .i_rd_waddr(rf_writeAddress),
      .i_rd_wen  (reg2_regWrite),
      .i_rd_wdata(WriteDataReg)
  );



/* 
 ID/EX Piepline Register
*/
  reg [31:0] reg1_PC_plus4;
  reg [31:0] reg1_current_PC;
  reg [31:0] reg0_immediate_val;
  reg [2:0] reg0_func3_val;
  reg reg0_branch_C;
  reg reg0_MemRead_C;
  reg [1:0] reg0_Data_sel_C;
  reg reg0_MemWrite_C;
  reg [31:0] reg0_ALU_operand1;
  reg [31:0] reg0_ALU_operand2;
  reg [31:0] reg0_Mem_WD;
  reg [2:0] reg0_ALUop_C;
  reg [3:0] reg0_func_val;
  reg [6:0] reg0_OP;
  reg reg1_retire_valid; 


reg [31:0] reg0_regData1;
reg [31:0] reg0_regData2;
  //include mux to control WB, M and EX inputs 

  always @(posedge i_clk) begin
    if (i_rst || Mux_sel || flush) begin
      reg1_current_PC    <= 32'd0;
      reg1_PC_plus4      <= 32'd0;
      reg0_immediate_val <= 32'd0;
      reg0_func3_val     <= 3'd0;
      reg0_jal_C         <= 1'd0;
      reg0_jalr_C        <= 1'd0;
      reg0_branch_C      <= 1'd0;
      reg0_regWrite      <= 1'd0;
      reg0_MemRead_C     <= 1'd0; 
      reg0_Data_sel_C    <= 2'd0; 
      reg0_MemWrite_C    <= 1'd0;
      reg0_ALU_operand1  <= 32'd0;
      reg0_ALU_operand2  <= 32'd0;
      reg0_Mem_WD        <= 32'd0;
      reg0_ALUop_C       <= 3'd0;
      reg0_func_val      <= 4'd0;
      reg0_OP            <= 7'd0;
      reg1_curr_instruct <= 32'd0;
      reg1_retire_valid  <= 1'd0;
      reg0_regData1      <= 32'd0;
      reg0_regData2      <=32'd0;

    end else begin
      reg1_current_PC    <= reg0_current_PC;
      reg1_PC_plus4      <= reg0_PC_plus4;
      reg0_immediate_val <= immediate_val;
      reg0_func3_val     <= func3_val;
      reg0_jal_C         <= jal_C;
      reg0_jalr_C        <= jalr_C;
      reg0_branch_C      <= branch_C;
      reg0_regWrite      <= regWrite;
      reg0_MemRead_C     <= MemRead_C;
      reg0_Data_sel_C    <= Data_sel_C;
      reg0_MemWrite_C    <= MemWrite_C;
      reg0_ALU_operand1  <= ALU_operand1;
      reg0_ALU_operand2  <= ALU_operand2;
      reg0_Mem_WD        <= Mem_WD;
      reg0_ALUop_C       <= ALUop_C;
      reg0_func_val      <= func_val;
      reg0_OP            <= reg0_curr_instruct[6:0];
      reg1_curr_instruct <= reg0_curr_instruct; 
      reg1_retire_valid  <= reg0_retire_valid;
      reg0_regData1      <= regData1;
      reg0_regData2      <= regData2;      
    end 
 end


  /* 
 Instantiate EX section of proccesor 
*/
  EX execute_I (
      .i_pc(reg1_current_PC),      //input- Current PC input should be added to immediate (used for branch instructions)
      .func3(reg0_func3_val),  //input- func 3 input for branch logic block (branch.v file)
      .i_jal(reg0_jal_C),  //input- control signal for branch logic block
      .i_jalr(reg0_jalr_C),  //input- control signal for branch logic block
      .i_branch(reg0_branch_C),  //input- control signal for branch logic block
      .i_ALUOp(reg0_ALUop_C),  //input- input to ALU CTRL unit
      .i_op1(reg0_ALU_operand1),  //input- ALU operand1
      .i_op2(reg0_ALU_operand2),  //input- ALU operand2
      .i_imm(reg0_immediate_val),        //input- i_imm is used for adding to current PC if we are in I instruction i_op2 will be input as immediate already
      .func(reg0_func_val),  //input- combination of func7 and func 3 used by ALU control

      .o_result(ALU_result),  //output- ALU result
      .o_PC_Select(PC_MUX_SEL),     //output- MUX select signals from branch logic unit used to select next PC
      .o_inc_pc(PC_offset)          //output- The current PC + Immediate (used for branch adress calculation)
  );

  
assign JB_PC = (PC_MUX_SEL[1]) ? PC_offset :  ALU_result;

wire byte_hw_unsigned;
wire [3:0] mask;
wire [31:0] WriteDataMem;
reg [3:0]  reg1_mask;
reg reg1_byte_hw_unsigned;

S_extend dataEXT(
  .i_mask(mask),         
  .i_unsign(byte_hw_unsigned),
  .i_old_mask(reg1_mask),
  .i_old_unsign(reg1_byte_hw_unsigned), 

  .i_Rs2Data(reg0_Mem_WD),                 //register data input 
  .o_Memdata(WriteDataMem),           //aligned output based on mask 

  .i_WB(WB_DATA),
  .o_regData(WriteDataReg)
);


wire [31:0] aligned_address;
  mask_gen mask_gen (
      .address(ALU_result),
      .func3(reg0_func3_val),
      .aligned_address(aligned_address),
      .o_unsigned(byte_hw_unsigned),
      .mask(mask),
      .opcode(reg0_OP)
  );


  /*
  EX/MEM Pipeline Register
  */
  reg [31:0] reg2_PC_plus4;
  reg [31:0] reg0_alu_result;
  reg [31:0] reg0_aligned_address; 
  reg [3:0] reg0_mask;
  reg reg0_byte_hw_unsigned;
  reg [31:0] reg0_ALU_result;
  reg [31:0] reg1_immediate_val; 
  reg reg1_MemRead_C;
  reg [1:0] reg1_Data_sel_C; 
  reg reg1_MemWrite_C; 
  reg [31:0] reg0_WriteDataMem; 
  reg reg2_retire_valid;
  reg [31:0] reg2_current_PC;

  reg [31:0] reg1_regData1;
  reg [31:0] reg1_regData2;

  always @(posedge i_clk) begin
    if (i_rst) begin
      reg1_jal_C<=1'b0;
      reg2_PC_plus4 <= 32'b0;
      reg0_aligned_address <= 32'b0;
      reg0_mask <= 4'b0;
      reg0_byte_hw_unsigned <= 1'b0;
      reg0_ALU_result <= 32'b0;
      reg1_immediate_val <= 32'd0;
      reg1_regWrite <= 1'd0;
      reg1_MemRead_C <= 1'd0;
      reg1_Data_sel_C <= 2'd0;
      reg1_MemWrite_C <= 1'd0;
      reg0_WriteDataMem <= 32'd0;
      reg2_curr_instruct <= 32'd0;
      reg2_retire_valid  <= 1'd0;
      reg2_current_PC    <= 32'd0;
      reg1_regData2     <= 32'd0;
      reg1_regData1     <= 32'd0;   

    end else begin
      reg1_jal_C<=reg0_jal_C;
      reg2_PC_plus4 <= reg1_PC_plus4;
      reg0_aligned_address <= aligned_address;
      reg0_mask <= mask;
      reg0_byte_hw_unsigned <= byte_hw_unsigned;
      reg0_ALU_result <= ALU_result;
      reg1_immediate_val <= reg0_immediate_val;
      reg1_regWrite <= reg0_regWrite;
      reg1_MemRead_C <= reg0_MemRead_C;
      reg1_Data_sel_C <= reg0_Data_sel_C;
      reg1_MemWrite_C <= reg0_MemWrite_C;
      reg0_WriteDataMem <= WriteDataMem;
      reg2_curr_instruct <= reg1_curr_instruct;
      reg2_retire_valid  <= reg1_retire_valid;
      reg2_current_PC    <= reg1_current_PC;
      reg1_regData2     <= reg0_regData2;
      reg1_regData1     <= reg0_regData1;       
    end
  end

  /* 
 Instantiate MEM section of proccesor  (actual memory access done outside MEM module)
*/




  assign o_dmem_addr = reg0_aligned_address;  //assign memory adress port to ALU result  
  assign o_dmem_ren  = reg1_MemRead_C;   //assign Memory Read enable signal 
  assign o_dmem_wen  = reg1_MemWrite_C;  //assign Memory Write enable signal 
  assign o_dmem_wdata = reg0_WriteDataMem;     //assign Memory Write data port to register output #2
  assign MEM_DATA = i_dmem_rdata;    //data returned from memory 



/* 
 MEM/WB pipeline register  
*/
reg [1:0]  reg2_Data_sel_C;
reg [31:0] reg0_MEM_DATA;
reg [31:0] reg1_ALU_result;
reg [31:0] reg2_immediate_val;
reg [31:0] reg3_PC_plus4; 
reg reg3_retire_valid;
reg [31:0] reg3_current_PC;
reg [31:0] reg1_aligned_address;
reg reg2_MemRead_C;
reg reg2_MemWrite_C;
reg [31:0] reg1_WriteDataMem;

reg [31:0] reg2_regData1;
reg [31:0] reg2_regData2;

always @(posedge i_clk) begin
    if (i_rst)begin
      reg2_regWrite         <= 1'd0;
      reg2_Data_sel_C       <= 2'd0;
      reg0_MEM_DATA         <= 32'd0; 
      reg1_ALU_result       <= 32'd0;
      reg2_immediate_val    <= 32'd0;
      reg3_PC_plus4         <= 32'd0;
      reg1_mask             <= 4'd0;
      reg1_byte_hw_unsigned <= 1'd0;
      reg3_curr_instruct    <= 32'd0; 
      reg3_retire_valid     <= 1'd0;
      reg3_current_PC       <= 32'd0;  
      reg1_aligned_address  <= 32'd0;
      reg2_MemRead_C        <= 1'd0; 
      reg2_MemWrite_C       <= 1'd0;
      reg1_WriteDataMem     <= 32'd0;
      reg2_regData1         <= 32'd0;
      reg2_regData2         <= 32'd0;   
    end else begin
      reg2_regWrite         <= reg1_regWrite;
      reg2_Data_sel_C       <= reg1_Data_sel_C; 
      reg0_MEM_DATA         <= MEM_DATA;
      reg1_ALU_result       <= reg0_ALU_result;
      reg2_immediate_val    <= reg1_immediate_val; 
      reg3_PC_plus4         <= reg2_PC_plus4;
      reg1_mask             <= reg0_mask;
      reg1_byte_hw_unsigned <= reg0_byte_hw_unsigned;
      reg3_curr_instruct    <= reg2_curr_instruct; 
      reg3_retire_valid     <= reg2_retire_valid;
      reg3_current_PC       <= reg2_current_PC;
      reg1_aligned_address  <= reg0_aligned_address;
      reg2_MemRead_C        <= reg1_MemRead_C;
      reg2_MemWrite_C       <= reg1_MemWrite_C;
      reg1_WriteDataMem     <= reg0_WriteDataMem; 
      reg2_regData1         <= reg1_regData1;
      reg2_regData2         <= reg1_regData2;
    end 
 end


  /* 
 Instantiate WB section of proccesor 
*/
  WB writeback (

      .i_MemData(MEM_DATA),  //input-  data coming from Memory
      .i_AluRslt(reg1_ALU_result),  //input- ALU operation result 
      .i_imm(reg2_immediate_val),  //input- output from immediate generator 
      .i_PC4(reg3_PC_plus4),  //input- incremented PC (used to save jump return adress in register)
      .i_MUXsel(reg2_Data_sel_C),  //input- MUX select signals coming from control unit 

      .o_dataSel(WB_DATA)        //output- data selected from mux to feedback into write port of Register file
  );


  /*
THIS section still needs to be checked and filled in properly (some values are being used as placeholders for now)
We can add extra output signals from modules to connect below 
*/
  assign o_dmem_mask = reg0_mask; //this used to control half word/byte loads and write (set to full word only for now)


  assign o_retire_valid = reg3_retire_valid &  ~i_rst; //one instruction should be done every cycle
  assign o_retire_inst = reg3_curr_instruct;
  assign o_retire_trap = 1'b0;  // implement trap detection later
  assign o_retire_halt = (reg3_curr_instruct == 32'h00100073);  // detect ebreak in ID stage 

  // retire register addresses (taken directly from the instruction fields)
  assign o_retire_rs1_raddr = reg3_curr_instruct[19:15];
  assign o_retire_rs2_raddr = reg3_curr_instruct[24:20];
  assign o_retire_rd_waddr = rf_writeAddress;

  // retire register read data 
  // Ideally use the raw register-file read data
  assign o_retire_rs1_rdata = reg2_regData1;
  assign o_retire_rs2_rdata = reg2_regData2;

  // retire write-back info (what is written back this cycle)
  assign o_retire_rd_wdata = WriteDataReg;

  // retire PC values
  assign o_retire_pc = reg3_current_PC;
  assign o_retire_next_pc = next_PC;

  assign o_retire_dmem_addr = reg1_aligned_address; 
  assign o_retire_dmem_ren = reg2_MemRead_C;
  assign o_retire_dmem_wen = reg2_MemWrite_C;
  assign o_retire_dmem_mask = reg1_mask; 
  assign o_retire_dmem_wdata = reg1_WriteDataMem; 
  assign o_retire_dmem_rdata = MEM_DATA; 


endmodule
`default_nettype wire
