module hazard();


endmodule